// hazard unit; checks current pipeline state for hazards
// and either stalls appropriately or forwards needed data
// by controlling forwarding muxes.
module hazard (
);

endmodule