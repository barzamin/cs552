module writeback (
    output wire err
);

    assign err = 1'b0;
endmodule
