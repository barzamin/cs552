module flop_mem2wb(
    input wire clk,
    input wire rst,
);

endmodule