module cache_fsm();

endmodule
