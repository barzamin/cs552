module flop_id2ex(
    input wire clk,
    input wire rst,
);

endmodule