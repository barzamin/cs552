module flop_if2id(
    input wire clk,
    input wire rst,
);

endmodule