module flop_ex2mem(
    input wire clk,
    input wire rst,
);

endmodule